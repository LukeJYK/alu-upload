-v200x -64bit -gui -access r
eecs361/lib/xor_gate.vhd
eecs361/lib/and_gate.vhd
eecs361/lib/or_gate.vhd
eecs361/lib/not_gate.vhd
eecs361/lib/xor_gate_32.vhd
eecs361/lib/mux.vhd
eecs361/lib/mux_n.vhd
eecs361/lib/eecs361_gates.vhd
eecs361/lib/eecs361.vhd
full_adder.vhd
half_adder.vhd
adder_32.vhd
sub_32.vhd
rshift.vhd
lshift.vhd
alu_32.vhd
mux_16.vhd
mux_16single.vhd
slt_32.vhd
sltu_32.vhd
zero_detect.vhd
alu_32_t.vhd
-top alu_32_t
