-v200x -64bit -gui -access r
eecs361/lib/xor_gate.vhd
eecs361/lib/and_gate.vhd
eecs361/lib/or_gate.vhd
eecs361/lib/eecs361_gates.vhd
full_adder.vhd 
half_adder.vhd
adder_8bit.vhd
adder_32bit.vhd
adder_32bit_t.vhd
-top adder_32bit_t

