-v200x -64bit -gui -access r
./eecs361/lib/eecs361_gates.vhd
half_adder.vhd
half_adder_t.vhd -top half_adder_t

