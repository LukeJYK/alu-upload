-v200x -64bit -gui -access r
eecs361/lib/xor_gate.vhd
eecs361/lib/and_gate.vhd
eecs361/lib/or_gate.vhd
eecs361/lib/xor_gate_32
eecs361/lib/mux
eecs361/lib/mux_n
eecs361/lib/eecs361_gates.vhd
eecs361/lib/eecs361.vhd
full_adder.vhd
half_adder.vhd
adder_8bit.vhd
adder_32bit.vhd
add_sub32bit.vhd
add_sub32bit_t.vhd
-top add_sub32bit_t
